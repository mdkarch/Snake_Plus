// sram.v

// Generated using ACDS version 12.1 177 at 2013.04.02.15:29:09

`timescale 1 ps / 1 ps
module sram (
		input  wire        chipselect, // avalon_slave_0.chipselect
		input  wire        write,      //               .write
		input  wire        read,       //               .read
		input  wire [17:0] address,    //               .address
		output wire [15:0] readdata,   //               .readdata
		input  wire [15:0] writedata,  //               .writedata
		input  wire [1:0]  byteenable, //               .byteenable
		inout  wire [15:0] SRAM_DQ,    //    conduit_end.export
		output wire [17:0] SRAM_ADDR,  //               .export
		output wire        SRAM_UB_N,  //               .export
		output wire        SRAM_LB_N,  //               .export
		output wire        SRAM_WE_N,  //               .export
		output wire        SRAM_CE_N,  //               .export
		output wire        SRAM_OE_N   //               .export
	);

	de2_sram_controller sram_inst (
		.chipselect (chipselect), // avalon_slave_0.chipselect
		.write      (write),      //               .write
		.read       (read),       //               .read
		.address    (address),    //               .address
		.readdata   (readdata),   //               .readdata
		.writedata  (writedata),  //               .writedata
		.byteenable (byteenable), //               .byteenable
		.SRAM_DQ    (SRAM_DQ),    //    conduit_end.export
		.SRAM_ADDR  (SRAM_ADDR),  //               .export
		.SRAM_UB_N  (SRAM_UB_N),  //               .export
		.SRAM_LB_N  (SRAM_LB_N),  //               .export
		.SRAM_WE_N  (SRAM_WE_N),  //               .export
		.SRAM_CE_N  (SRAM_CE_N),  //               .export
		.SRAM_OE_N  (SRAM_OE_N)   //               .export
	);

endmodule
