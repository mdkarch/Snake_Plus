// vga.v

// Generated using ACDS version 12.1 177 at 2013.04.03.11:55:04

`timescale 1 ps / 1 ps
module vga (
		input  wire        clk,        //          clock.clk
		input  wire        reset_n,    //          reset.reset_n
		input  wire        read,       // avalon_slave_0.read
		input  wire        write,      //               .write
		input  wire        chipselect, //               .chipselect
		input  wire [2:0]  address,    //               .address
		output wire [15:0] readdata,   //               .readdata
		input  wire [15:0] writedata,  //               .writedata
		output wire        VGA_CLK,    //    conduit_end.export
		output wire        VGA_HS,     //               .export
		output wire        VGA_VS,     //               .export
		output wire        VGA_BLANK,  //               .export
		output wire        VGA_SYNC,   //               .export
		output wire [9:0]  VGA_R,      //               .export
		output wire [9:0]  VGA_G,      //               .export
		output wire [9:0]  VGA_B,      //               .export
		output wire [15:0] leds        //               .export
	);

	snake_plus_vga vga_inst (
		.clk        (clk),        //          clock.clk
		.reset_n    (reset_n),    //          reset.reset_n
		.read       (read),       // avalon_slave_0.read
		.write      (write),      //               .write
		.chipselect (chipselect), //               .chipselect
		.address    (address),    //               .address
		.readdata   (readdata),   //               .readdata
		.writedata  (writedata),  //               .writedata
		.VGA_CLK    (VGA_CLK),    //    conduit_end.export
		.VGA_HS     (VGA_HS),     //               .export
		.VGA_VS     (VGA_VS),     //               .export
		.VGA_BLANK  (VGA_BLANK),  //               .export
		.VGA_SYNC   (VGA_SYNC),   //               .export
		.VGA_R      (VGA_R),      //               .export
		.VGA_G      (VGA_G),      //               .export
		.VGA_B      (VGA_B),      //               .export
		.leds       (leds)        //               .export
	);

endmodule
