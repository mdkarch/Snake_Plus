// de2_audio_0.v

// Generated using ACDS version 12.1 177 at 2013.04.22.12:05:10

`timescale 1 ps / 1 ps
module de2_audio_0 (
		input  wire        clk,         //          clock.clk
		input  wire        reset_n,     //          reset.reset_n
		input  wire        read,        // avalon_slave_0.read
		input  wire        write,       //               .write
		input  wire        chipselect,  //               .chipselect
		input  wire [2:0]  address,     //               .address
		output wire [15:0] readdata,    //               .readdata
		input  wire [15:0] writedata,   //               .writedata
		output wire        AUD_ADCLRCK, //    conduit_end.export
		input  wire        AUD_ADCDAT,  //               .export
		output wire        AUD_DACLRCK, //               .export
		output wire        AUD_DACDAT,  //               .export
		inout  wire        AUD_BCLK,    //               .export
		output wire        AUD_XCK,     //               .export
		input  wire        iCLK,        //               .export
		input  wire        iRST_N,      //               .export
		output wire        I2C_SCLK,    //               .export
		inout  wire        I2C_SDAT     //               .export
	);

	de2_audio de2_audio_0_inst (
		.clk         (clk),         //          clock.clk
		.reset_n     (reset_n),     //          reset.reset_n
		.read        (read),        // avalon_slave_0.read
		.write       (write),       //               .write
		.chipselect  (chipselect),  //               .chipselect
		.address     (address),     //               .address
		.readdata    (readdata),    //               .readdata
		.writedata   (writedata),   //               .writedata
		.AUD_ADCLRCK (AUD_ADCLRCK), //    conduit_end.export
		.AUD_ADCDAT  (AUD_ADCDAT),  //               .export
		.AUD_DACLRCK (AUD_DACLRCK), //               .export
		.AUD_DACDAT  (AUD_DACDAT),  //               .export
		.AUD_BCLK    (AUD_BCLK),    //               .export
		.AUD_XCK     (AUD_XCK),     //               .export
		.iCLK        (iCLK),        //               .export
		.iRST_N      (iRST_N),      //               .export
		.I2C_SCLK    (I2C_SCLK),    //               .export
		.I2C_SDAT    (I2C_SDAT)     //               .export
	);

endmodule
