library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package sounds is

	type sound1_type is array(0 to 4106) of unsigned(15 downto 0);
	type sound2_type is array(0 to 1366) of unsigned(15 downto 0);
	
	
	constant sound1 : sound1_type :=	 (
		X"0000", X"1172", X"102F", X"0F02", X"0DEC", X"0CE9", 
		X"E999", X"EB39", X"ECBB", X"EE21", X"EF6D", X"F0A1", 
		X"F1BF", X"14BC", X"133A", X"11D5", X"108A", X"0F57", 
		X"EACA", X"EC55", X"EDC2", X"EF15", X"F04F", X"F173", 
		X"F281", X"1506", X"137F", X"1215", X"10C5", X"0F8E", 
		X"EB19", X"EC9D", X"EE06", X"EF54", X"F089", X"F1A9", 
		X"0A21", X"14E3", X"135F", X"11F8", X"10AA", X"0F74", 
		X"EB5C", X"ECDC", X"EE3F", X"EF89", X"F0BB", X"F1D7", 
		X"163A", X"149D", X"131E", X"11BB", X"1072", X"0F40", 
		X"EBB3", X"ED2C", X"EE8A", X"EFCE", X"F0FB", X"F212", 
		X"15C2", X"142E", X"12B7", X"115B", X"1019", X"F449", 
		X"EC29", X"ED9A", X"EEEF", X"F02C", X"F153", X"F263", 
		X"1536", X"13AC", X"123F", X"10EC", X"0FB2", X"EB33", 
		X"ECB5", X"EE1C", X"EF68", X"F09C", X"F1BA", X"126F", 
		X"1495", X"1317", X"11B4", X"106C", X"0F3B", X"EBDF", 
		X"ED55", X"EEAF", X"EFF1", X"F11B", X"F230", X"1570", 
		X"13E1", X"1270", X"111A", X"0FDC", X"EB18", X"EC9C", 
		X"EE04", X"EF52", X"F088", X"F1A8", X"0D72", X"149B", 
		X"131D", X"11BA", X"1070", X"0F3F", X"EBF5", X"ED69", 
		X"EEC3", X"F003", X"F12C", X"F23F", X"1531", X"13A8", 
		X"123B", X"10E8", X"0FAE", X"EB6B", X"ECEA", X"EE4C", 
		X"EF95", X"F0C6", X"F1E1", X"15B5", X"1422", X"12AC", 
		X"1151", X"100F", X"EEFE", X"EC80", X"EDEA", X"EF3A", 
		X"F072", X"F193", X"09AC", X"1487", X"130A", X"11A8", 
		X"1060", X"0F30", X"EC2C", X"ED9C", X"EEF2", X"F02F", 
		X"F155", X"F265", X"14D5", X"1352", X"11EB", X"109E", 
		X"0F69", X"EBEF", X"ED64", X"EEBD", X"EFFE", X"F127", 
		X"F23B", X"150A", X"1383", X"1219", X"10C9", X"0F91", 
		X"EBC9", X"ED41", X"EE9D", X"EFE0", X"F10C", X"F222", 
		X"1527", X"139E", X"1231", X"10E0", X"0FA6", X"EBBC", 
		X"ED35", X"EE92", X"EFD6", X"F102", X"F219", X"152A", 
		X"13A1", X"1234", X"10E2", X"0FA8", X"EBC7", X"ED3F", 
		X"EE9C", X"EFDF", X"F10A", X"F220", X"1514", X"138C", 
		X"1221", X"10D0", X"0F98", X"EBEB", X"ED60", X"EEBA", 
		X"EFFB", X"F125", X"F239", X"14E4", X"1360", X"11F8", 
		X"10AA", X"0F75", X"EC26", X"ED97", X"EEED", X"F02A", 
		X"F151", X"F261", X"149C", X"131E", X"11BA", X"1071", 
		X"0F40", X"EC78", X"EDE3", X"EF34", X"F06C", X"F18D", 
		X"0957", X"143D", X"12C5", X"1168", X"1025", X"EF67", 
		X"ECE0", X"EE44", X"EF8D", X"F0BF", X"F1DA", X"1554", 
		X"13C8", X"1258", X"1103", X"0FC7", X"EBD5", X"ED4C", 
		X"EEA7", X"EFEA", X"F115", X"F22A", X"14B8", X"1338", 
		X"11D3", X"1088", X"0F54", X"EC6D", X"EDD9", X"EF2A", 
		X"F063", X"F185", X"092E", X"141F", X"12A9", X"114E", 
		X"100D", X"EB95", X"ED10", X"EE70", X"EFB6", X"F0E5", 
		X"F1FD", X"14F5", X"1370", X"1207", X"10B8", X"0F81", 
		X"EC55", X"EDC3", X"EF15", X"F050", X"F173", X"F5E9", 
		X"1426", X"12AF", X"1154", X"1012", X"EBAC", X"ED25", 
		X"EE84", X"EFC8", X"F0F6", X"F20D", X"14C9", X"1347", 
		X"11E1", X"1095", X"0F61", X"EC9A", X"EE03", X"EF51", 
		X"F087", X"F1A6", X"1396", X"13CC", X"125C", X"1107", 
		X"0FCB", X"EC11", X"ED83", X"EEDB", X"F019", X"F141", 
		X"F253", X"1445", X"12CD", X"1170", X"102C", X"F22C", 
		X"ED1C", X"EE7B", X"EFC0", X"F0EE", X"F206", X"14AB", 
		X"132B", X"11C7", X"107D", X"0F4A", X"ECCA", X"EE2F", 
		X"EF7A", X"F0AD", X"F1CA", X"14F9", X"1374", X"120A", 
		X"10BB", X"0F85", X"EC8F", X"EDF9", X"EF48", X"F07E", 
		X"F19E", X"136E", X"13A6", X"1239", X"10E7", X"0FAD", 
		X"EC59", X"EDC6", X"EF19", X"F053", X"F176", X"08C0", 
		X"13CB", X"125B", X"1106", X"0FCA", X"EC3F", X"EDAE", 
		X"EF03", X"F03E", X"F163", X"F5BE", X"13D9", X"1269", 
		X"1113", X"0FD5", X"EC3E", X"EDAD", X"EF02", X"F03E", 
		X"F162", X"F5BA", X"13D0", X"1260", X"110B", X"0FCE", 
		X"EC55", X"EDC3", X"EF15", X"F050", X"F173", X"FBA9", 
		X"13C0", X"1251", X"10FD", X"0FC1", X"EC68", X"EDD4", 
		X"EF26", X"F05F", X"F181", X"0F17", X"138E", X"1223", 
		X"10D2", X"0F99", X"EC9F", X"EE07", X"EF55", X"F08B", 
		X"F1AA", X"14CC", X"134A", X"11E4", X"1097", X"0F63", 
		X"ECEE", X"EE51", X"EF99", X"F0CA", X"F1E5", X"147D", 
		X"1300", X"119F", X"1058", X"0C70", X"ED4B", X"EEA6", 
		X"EFE9", X"F114", X"F229", X"1413", X"129E", X"1144", 
		X"1004", X"EC39", X"EDA9", X"EEFE", X"F03A", X"F15F", 
		X"F5A6", X"139D", X"1230", X"10DE", X"0FA5", X"ECB9", 
		X"EE1F", X"EF6B", X"F09F", X"F1BD", X"1491", X"1313", 
		X"11B1", X"1068", X"0F38", X"ED4D", X"EEA8", X"EFEA", 
		X"F115", X"F22A", X"13FA", X"1287", X"112F", X"0FF0", 
		X"EC6D", X"EDD8", X"EF2A", X"F063", X"F185", X"1113", 
		X"1346", X"11E0", X"1094", X"0F60", X"ED22", X"EE81", 
		X"EFC6", X"F0F3", X"F20B", X"140A", X"1296", X"113D", 
		X"0FFD", X"EC75", X"EDE0", X"EF31", X"F069", X"F18B", 
		X"1107", X"1339", X"11D4", X"1089", X"0F56", X"ED3E", 
		X"EE9B", X"EFDE", X"F10A", X"F220", X"13D3", X"1263", 
		X"110D", X"0FD1", X"ECB3", X"EE19", X"EF66", X"F09A", 
		X"F1B8", X"145B", X"12E1", X"1182", X"103D", X"FC5F", 
		X"EDAB", X"EF00", X"F03C", X"F161", X"F594", X"135C", 
		X"11F4", X"10A7", X"0F71", X"ED48", X"EEA4", X"EFE6", 
		X"F112", X"F227", X"13BE", X"1250", X"10FB", X"0FC0", 
		X"ECE6", X"EE49", X"EF92", X"F0C4", X"F1DF", X"1413", 
		X"129E", X"1144", X"1004", X"EC9E", X"EE07", X"EF55", 
		X"F08A", X"F1AA", X"1464", X"12E9", X"118A", X"1044", 
		X"08E3", X"EDC0", X"EF13", X"F04E", X"F172", X"0BCE", 
		X"1314", X"11B2", X"1069", X"0F38", X"ED9B", X"EEF1", 
		X"F02E", X"F154", X"F265", X"133D", X"11D8", X"108C", 
		X"0F59", X"ED86", X"EEDD", X"F01C", X"F143", X"F255", 
		X"134D", X"11E6", X"109A", X"0F65", X"ED74", X"EECD", 
		X"F00C", X"F135", X"F248", X"134E", X"11E7", X"109B", 
		X"0F66", X"ED7D", X"EED5", X"F014", X"F13C", X"F24E", 
		X"134A", X"11E3", X"1097", X"0F63", X"ED95", X"EEEB", 
		X"F028", X"F14F", X"F260", X"132B", X"11C7", X"107D", 
		X"0F4A", X"EDAF", X"EF04", X"F03F", X"F164", X"FA65", 
		X"12FE", X"119D", X"1056", X"0F26", X"EDD3", X"EF25", 
		X"F05E", X"F181", X"108E", X"12C5", X"1168", X"1025", 
		X"F68D", X"EE12", X"EF5F", X"F094", X"F1B3", X"13FC", 
		X"1289", X"1130", X"0FF1", X"ECFD", X"EE5E", X"EFA6", 
		X"F0D6", X"F1F0", X"13A1", X"1234", X"10E2", X"0FA8", 
		X"ED51", X"EEAC", X"EFEE", X"F119", X"F22E", X"1338", 
		X"11D3", X"1088", X"0F55", X"EDBE", X"EF12", X"F04C", 
		X"F170", X"0781", X"12CD", X"1170", X"102C", X"F6C2", 
		X"EE37", X"EF82", X"F0B4", X"F1D1", X"13BA", X"124B", 
		X"10F7", X"0FBC", X"ED55", X"EEB0", X"EFF2", X"F11C", 
		X"F231", X"1322", X"11BF", X"1075", X"0F43", X"EDEE", 
		X"EF3E", X"F075", X"F196", X"1245", X"128B", X"1132", 
		X"0FF3", X"ED21", X"EE7F", X"EFC5", X"F0F2", X"F20A", 
		X"134E", X"11E7", X"109B", X"0F66", X"EDD1", X"EF23", 
		X"F05D", X"F17F", X"0B5B", X"129F", X"1145", X"1004", 
		X"EEF2", X"EE79", X"EFBF", X"F0ED", X"F205", X"133B", 
		X"11D6", X"108B", X"0F57", X"EDE9", X"EF39", X"F071", 
		X"F192", X"1223", X"126A", X"1114", X"0FD7", X"ED54", 
		X"EEAF", X"EFF1", X"F11B", X"F230", X"12F3", X"1193", 
		X"104C", X"0F1D", X"EE38", X"EF83", X"F0B5", X"F1D1", 
		X"137A", X"1210", X"10C0", X"0F89", X"EDCE", X"EF20", 
		X"F059", X"F17C", X"0732", X"1287", X"112F", X"0FF0", 
		X"ED5B", X"EEB5", X"EFF7", X"F121", X"F235", X"12EF", 
		X"118F", X"1049", X"0F1A", X"EE60", X"EFA7", X"F0D7", 
		X"F1F1", X"1353", X"11EC", X"109F", X"0F6A", X"EE05", 
		X"EF53", X"F089", X"F1A9", X"1396", X"122A", X"10D9", 
		X"0FA0", X"EDCA", X"EF1D", X"F056", X"F17A", X"0703", 
		X"1268", X"1112", X"0FD5", X"ED8D", X"EEE4", X"F022", 
		X"F149", X"F25B", X"1296", X"113C", X"0FFC", X"F14A", 
		X"EEB3", X"EFF4", X"F11E", X"F233", X"12B7", X"115B", 
		X"1019", X"0268", X"EE9B", X"EFDE", X"F10A", X"F220", 
		X"12D5", X"1177", X"1033", X"0F06", X"EE81", X"EFC6", 
		X"F0F4", X"F20C", X"12E2", X"1183", X"103E", X"0F10", 
		X"EE7F", X"EFC5", X"F0F2", X"F20A", X"12EA", X"118A", 
		X"1045", X"0F16", X"EE8C", X"EFD0", X"F0FD", X"F214", 
		X"12E8", X"1189", X"1043", X"0F15", X"EE93", X"EFD7", 
		X"F103", X"F21A", X"12D3", X"1176", X"1031", X"0C98", 
		X"EEB1", X"EFF2", X"F11D", X"F232", X"12B9", X"115E", 
		X"101B", X"032D", X"EECC", X"F00B", X"F134", X"F247", 
		X"128E", X"1135", X"0FF6", X"EF7E", X"EEFE", X"F03A", 
		X"F15F", X"F26F", X"125E", X"1109", X"0FCC", X"EDDB", 
		X"EF2C", X"F065", X"F187", X"06AC", X"121E", X"10CD", 
		X"0F95", X"EE14", X"EF61", X"F096", X"F1B4", X"1337", 
		X"11D2", X"1087", X"0F54", X"EE67", X"EFAE", X"F0DD", 
		X"F1F6", X"12E3", X"1184", X"103E", X"0F11", X"EEB6", 
		X"EFF7", X"F121", X"F236", X"127F", X"1127", X"0FE8", 
		X"EF9C", X"EF1B", X"F055", X"F178", X"F551", X"1218", 
		X"10C8", X"0F90", X"EE31", X"EF7C", X"F0AF", X"F1CB", 
		X"1305", X"11A3", X"105C", X"0F2C", X"EEAE", X"EFF0", 
		X"F11A", X"F22F", X"1285", X"112D", X"0FEE", X"F1C1", 
		X"EF25", X"F05E", X"F181", X"F978", X"11F8", X"10AA", 
		X"0F74", X"EE69", X"EFB0", X"F0DF", X"F1F8", X"12C7", 
		X"116A", X"1026", X"0EFA", X"EEF6", X"F033", X"F159", 
		X"F269", X"1222", X"10D1", X"0F98", X"EE4D", X"EF96", 
		X"F0C7", X"F1E2", X"12DC", X"117D", X"1038", X"0F0B", 
		X"EEF0", X"F02D", X"F153", X"F264", X"1220", X"10CF", 
		X"0F97", X"EE4A", X"EF94", X"F0C5", X"F1E0", X"12BB", 
		X"115F", X"101C", X"0EF1", X"EEFD", X"F03A", X"F15F", 
		X"F26F", X"11E9", X"109C", X"0F67", X"EE7D", X"EFC3", 
		X"F0F1", X"F208", X"1273", X"111C", X"0FDE", X"F46C", 
		X"EF47", X"F07E", X"F19E", X"0F56", X"1191", X"104A", 
		X"0F1C", X"EEDF", X"F01D", X"F144", X"F256", X"1204", 
		X"10B5", X"0F7E", X"EE72", X"EFB8", X"F0E7", X"F1FF", 
		X"1278", X"1121", X"0FE3", X"F48B", X"EF60", X"F095", 
		X"F1B4", X"0F52", X"1188", X"1042", X"0F14", X"EF01", 
		X"F03D", X"F162", X"F272", X"11DF", X"1093", X"0F5F", 
		X"EEB7", X"EFF9", X"F123", X"F237", X"1233", X"10E1", 
		X"0FA8", X"EE69", X"EFB0", X"F0DF", X"F1F9", X"1277", 
		X"1120", X"0FE2", X"F820", X"EF6D", X"F0A1", X"F1BF", 
		X"12AF", X"1154", X"1012", X"0EE7", X"EF42", X"F079", 
		X"F19A", X"05DD", X"1185", X"103F", X"0F11", X"EF14", 
		X"F04F", X"F173", X"F281", X"11B6", X"106D", X"0F3B", 
		X"EEE6", X"F024", X"F14B", X"F25C", X"11D7", X"108B", 
		X"0F58", X"EECF", X"F00F", X"F137", X"F24A", X"11F4", 
		X"10A7", X"0F71", X"EEB6", X"EFF7", X"F121", X"F236", 
		X"1201", X"10B2", X"0F7C", X"EEA3", X"EFE5", X"F111", 
		X"F226", X"1200", X"10B2", X"0F7B", X"EEAA", X"EFEC", 
		X"F117", X"F22C", X"11FD", X"10AE", X"0F78", X"EEB0", 
		X"EFF1", X"F11C", X"F231", X"11F8", X"10AA", X"0F75", 
		X"EEC6", X"F006", X"F12F", X"F242", X"11EC", X"109F", 
		X"0F6A", X"EED7", X"F016", X"F13E", X"F250", X"11CE", 
		X"1083", X"0F50", X"EEEE", X"F02B", X"F151", X"F262", 
		X"11A3", X"105B", X"0F2B", X"EF1E", X"F058", X"F17B", 
		X"F289", X"1175", X"1031", X"0F04", X"EF4C", X"F082", 
		X"F1A2", X"F90B", X"1147", X"1006", X"0EDC", X"EF89", 
		X"F0BB", X"F1D7", X"10BF", X"1112", X"0FD5", X"04C1", 
		X"EFC1", X"F0EF", X"F207", X"121D", X"10CD", X"0F94", 
		X"EEBC", X"EFFD", X"F127", X"F23B", X"11C6", X"107C", 
		X"0F4A", X"EF05", X"F041", X"F165", X"F275", X"1175", 
		X"1031", X"0F04", X"EF60", X"F095", X"F1B4", X"055E", 
		X"1120", X"0FE2", X"0EBA", X"EFB5", X"F0E4", X"F1FD", 
		X"120B", X"10BC", X"0F85", X"EECF", X"F00F", X"F137", 
		X"F24A", X"1194", X"104D", X"0F1E", X"EF47", X"F07D", 
		X"F19E", X"F2A9", X"112D", X"0FEE", X"0EC6", X"EFB3", 
		X"F0E2", X"F1FB", X"1204", X"10B5", X"0F7F", X"EEE2", 
		X"F020", X"F147", X"F259", X"1179", X"1034", X"0F07", 
		X"EF6D", X"F0A1", X"F1BF", X"09A9", X"10EF", X"0FB4", 
		X"04D5", X"EFF2", X"F11C", X"F231", X"11B1", X"1069", 
		X"0F38", X"EF4C", X"F082", X"F1A2", X"F2AD", X"111E", 
		X"0FE0", X"0EB9", X"EFDD", X"F109", X"F21F", X"11C8", 
		X"107E", X"0F4B", X"EF36", X"F06E", X"F18F", X"F29C", 
		X"1124", X"0FE6", X"0EBE", X"EFDF", X"F10B", X"F221", 
		X"11CB", X"1081", X"0F4E", X"EF47", X"F07E", X"F19E", 
		X"F2A9", X"1110", X"0FD3", X"0EAD", X"EFF0", X"F11B", 
		X"F230", X"11A7", X"105F", X"0F2F", X"EF71", X"F0A5", 
		X"F1C2", X"F550", X"10EA", X"0FB0", X"0528", X"F027", 
		X"F14E", X"F25F", X"1168", X"1025", X"0EF9", X"EFAA", 
		X"F0DA", X"F1F4", X"11DC", X"1090", X"0F5D", X"EF32", 
		X"F06B", X"F18C", X"F299", X"1103", X"0FC7", X"0EA2", 
		X"F00B", X"F134", X"F247", X"1174", X"1030", X"0F03", 
		X"EFA6", X"F0D6", X"F1F0", X"1032", X"108A", X"0F57", 
		X"EF44", X"F07B", X"F19C", X"F2A7", X"10E9", X"0FAF", 
		X"0E8B", X"F020", X"F147", X"F258", X"113C", X"0FFB", 
		X"0ED2", X"EFD9", X"F106", X"F21C", X"119D", X"1055", 
		X"0F26", X"EF8A", X"F0BC", X"F1D8", X"04AE", X"109E", 
		X"0F69", X"F0FF", X"F074", X"F195", X"F2A1", X"10DA", 
		X"0FA1", X"0C5A", X"F042", X"F166", X"F276", X"1124", 
		X"0FE5", X"0EBE", X"F007", X"F130", X"F243", X"115B", 
		X"1019", X"0EED", X"EFCF", X"F0FC", X"F213", X"1185", 
		X"103F", X"0F11", X"EFAF", X"F0DE", X"F1F8", X"0C0F", 
		X"1073", X"0F41", X"EF86", X"F0B8", X"F1D5", X"F54E", 
		X"1094", X"0F60", X"F123", X"F096", X"F1B4", X"F2BE", 
		X"10A7", X"0F72", X"F5AD", X"F089", X"F1A9", X"F2B4", 
		X"10C8", X"0F90", X"09A5", X"F076", X"F197", X"F2A3", 
		X"10D5", X"0F9C", X"0E7A", X"F065", X"F187", X"F294", 
		X"10E4", X"0FAA", X"0E87", X"F056", X"F179", X"F287", 
		X"10E4", X"0FAB", X"0E87", X"F04C", X"F170", X"F27F", 
		X"10D9", X"0FA0", X"0E7D", X"F05C", X"F17F", X"F28C", 
		X"10DB", X"0FA2", X"0E7F", X"F064", X"F186", X"F293", 
		X"10CA", X"0F92", X"0E70", X"F06F", X"F191", X"F29D", 
		X"10BA", X"0F83", X"0C4B", X"F08C", X"F1AB", X"F2B6", 
		X"10A5", X"0F70", X"0574", X"F0A5", X"F1C2", X"F2CB", 
		X"108E", X"0F5A", X"F5DD", X"F0BC", X"F1D8", X"F2DF", 
		X"1067", X"0F37", X"EFA8", X"F0D8", X"F1F2", X"0407", 
		X"1035", X"0F08", X"EFE0", X"F10B", X"F221", X"0FB5", 
		X"1010", X"0EE6", X"F00F", X"F137", X"F24A", X"1117", 
		X"0FD9", X"0EB3", X"F041", X"F165", X"F275", X"10DF", 
		X"0FA5", X"0E82", X"F083", X"F1A3", X"F2AE", X"10A1", 
		X"0F6C", X"09A2", X"F0C1", X"F1DC", X"F2E3", X"1063", 
		X"0F32", X"EFCF", X"F0FC", X"F214", X"08E7", X"1015", 
		X"0EEA", X"F014", X"F13C", X"F24F", X"10F9", X"0FBE", 
		X"0E99", X"F06F", X"F191", X"F29D", X"10AA", X"0F75", 
		X"0E55", X"F0C2", X"F1DD", X"F2E4", X"104A", X"0F1B", 
		X"EFEB", X"F116", X"F22B", X"0DBE", X"0FEE", X"0EC5", 
		X"F044", X"F169", X"F278", X"10BD", X"0F85", X"0E65", 
		X"F0A2", X"F1C0", X"F2C9", X"1052", X"0F23", X"F19F", 
		X"F110", X"F225", X"0B8B", X"0FE7", X"0EBF", X"F054", 
		X"F177", X"F285", X"10B2", X"0F7C", X"0E5C", X"F0BF", 
		X"F1DB", X"F2E2", X"1032", X"0F05", X"F003", X"F12C", 
		X"F240", X"10F4", X"0FB9", X"0E94", X"F088", X"F1A8", 
		X"F2B2", X"1070", X"0F3E", X"05A8", X"F105", X"F21C", 
		X"F8A8", X"0FEE", X"0EC6", X"F05B", X"F17E", X"F28B", 
		X"1096", X"0F62", X"0E44", X"F0DD", X"F1F7", X"F2FC", 
		X"1006", X"0EDD", X"F048", X"F16D", X"F27C", X"10AD", 
		X"0F77", X"0E58", X"F0DA", X"F1F4", X"F2F9", X"1016", 
		X"0EEB", X"F040", X"F165", X"F275", X"10AB", X"0F75", 
		X"0E56", X"F0D6", X"F1F0", X"F2F5", X"1008", X"0EDE", 
		X"F054", X"F177", X"F286", X"109A", X"0F66", X"0E47", 
		X"F0F7", X"F20F", X"F312", X"0FF1", X"0EC8", X"F072", 
		X"F193", X"F29F", X"1071", X"0F3F", X"0E24", X"F118", 
		X"F22D", X"F89B", X"0FBC", X"0E98", X"F0AA", X"F1C7", 
		X"F2D0", X"1039", X"0F0B", X"F3F1", X"F15C", X"F26C", 
		X"10B7", X"0F80", X"0E60", X"F0EC", X"F204", X"F308", 
		X"0FE9", X"0EC2", X"F07E", X"F19E", X"F2AA", X"1058", 
		X"0F28", X"0C12", X"F137", X"F24A", X"0B30", X"0F85", 
		X"0E64", X"F0D3", X"F1ED", X"F2F3", X"0FE6", X"0EBF", 
		X"F06F", X"F190", X"F29D", X"103D", X"0F0F", X"097D", 
		X"F147", X"F259", X"0D42", X"0F6E", X"0E4F", X"F0F6", 
		X"F20D", X"F311", X"0FBC", X"0E97", X"F0A5", X"F1C3", 
		X"F2CB", X"100D", X"0EE3", X"F404", X"F177", X"F286", 
		X"1052", X"0F22", X"0E09", X"F140", X"F252", X"084D", 
		X"0F6F", X"0E50", X"F100", X"F217", X"F31A", X"0FB9", 
		X"0E95", X"F0BD", X"F1D9", X"F2E0", X"0FF4", X"0ECB", 
		X"F07D", X"F19E", X"F2A9", X"1032", X"0F05", X"0987", 
		X"F172", X"F281", X"106D", X"0F3B", X"0E20", X"F143", 
		X"F255", X"F89B", X"0F70", X"0E51", X"F112", X"F228", 
		X"F329", X"0F97", X"0E75", X"F0E5", X"F1FE", X"F303", 
		X"0FC0", X"0E9B", X"F0BA", X"F1D6", X"F2DD", X"0FDC", 
		X"0EB5", X"F0A4", X"F1C2", X"F2CB", X"1006", X"0EDC", 
		X"F6B6", X"F1A7", X"F2B2", X"102B", X"0EFF", X"0BF9", 
		X"F18A", X"F297", X"1041", X"0F13", X"0DFA", X"F171", 
		X"F27F", X"0D01", X"0F29", X"0E0F", X"F159", X"F269", 
		X"0813", X"0F31", X"0E17", X"F156", X"F266", X"F895", 
		X"0F47", X"0E2A", X"F14C", X"F25E", X"F58E", X"0F4A", 
		X"0E2D", X"F145", X"F257", X"F355", X"0F4E", X"0E32", 
		X"F13F", X"F252", X"F350", X"0F53", X"0E36", X"F14A", 
		X"F25B", X"F359", X"0F53", X"0E36", X"F150", X"F261", 
		X"F35F", X"0F51", X"0E35", X"F155", X"F266", X"F363", 
		X"0F40", X"0E24", X"F15E", X"F26E", X"F599", X"0F31", 
		X"0E17", X"F169", X"F278", X"F894", X"0F24", X"0E0A", 
		X"F175", X"F283", X"07F5", X"0F08", X"0DF1", X"F186", 
		X"F293", X"0CCA", X"0EF0", X"0DDA", X"F199", X"F2A5", 
		X"0FF4", X"0ECB", X"0BD1", X"F1C1", X"F2CA", X"0FDA", 
		X"0EB3", X"FAB1", X"F1E3", X"F2E9", X"0FBD", X"0E98", 
		X"F295", X"F202", X"F306", X"0F8F", X"0E6E", X"F10E", 
		X"F224", X"F326", X"0F64", X"0E46", X"F134", X"F247", 
		X"F346", X"0F2C", X"0E12", X"F16F", X"F27E", X"F59E", 
		X"0F02", X"0DEB", X"F1A3", X"F2AE", X"0CB3", X"0ED4", 
		X"0DC0", X"F1D4", X"F2DC", X"0FBC", X"0E98", X"F706", 
		X"F207", X"F30B", X"0F7E", X"0E5E", X"F128", X"F23C", 
		X"F33C", X"0F33", X"0E19", X"F174", X"F283", X"F37E", 
		X"0EF7", X"0DE0", X"F1BA", X"F2C3", X"0E57", X"0EB7", 
		X"0BC8", X"F1FB", X"F300", X"0F8B", X"0E6A", X"F12B", 
		X"F23F", X"F33F", X"0F3B", X"0E20", X"F174", X"F283", 
		X"F37E", X"0EEE", X"0DD8", X"F1CC", X"F2D4", X"0FC3", 
		X"0E9E", X"060B", X"F21E", X"F321", X"0F6C", X"0E4E", 
		X"F15D", X"F26D", X"F36A", X"0F08", X"0DF1", X"F1B5", 
		X"F2BF", X"0A71", X"0EA9", X"0D99", X"F20C", X"F30F", 
		X"0F6C", X"0E4D", X"F150", X"F262", X"F35F", X"0EFE", 
		X"0DE7", X"F1BF", X"F2C8", X"0A6A", X"0E9F", X"0BB7", 
		X"F225", X"F327", X"0F5C", X"0E3F", X"F177", X"F285", 
		X"F380", X"0EE7", X"0DD2", X"F1DF", X"F2E6", X"0F9A", 
		X"0E78", X"FB19", X"F246", X"F346", X"0F26", X"0E0C", 
		X"F19F", X"F2AB", X"F5B8", X"0EA8", X"0D97", X"F20E", 
		X"F311", X"0F4D", X"0E31", X"F16C", X"F27B", X"F376", 
		X"0ED2", X"0DBF", X"F1EE", X"F2F4", X"0F77", X"0E57", 
		X"F4EA", X"F269", X"F366", X"0EF5", X"0DDE", X"F1D7", 
		X"F2DE", X"0A46", X"0E76", X"0953", X"F250", X"F34F", 
		X"0F04", X"0DED", X"F1C1", X"F2CA", X"0044", X"0E79", 
		X"0D6C", X"F241", X"F341", X"0F0C", X"0DF4", X"F1C3", 
		X"F2CC", X"F893", X"0E7E", X"0D70", X"F250", X"F34F", 
		X"0F0A", X"0DF3", X"F1CE", X"F2D6", X"F89D", X"0E79", 
		X"0D6C", X"F259", X"F357", X"0EF6", X"0DE0", X"F1DB", 
		X"F2E2", X"0766", X"0E5A", X"0941", X"F26B", X"F367", 
		X"0ED9", X"0DC5", X"F1FF", X"F304", X"0DDA", X"0E3C", 
		X"F51A", X"F29A", X"F393", X"0EB4", X"0DA3", X"F22C", 
		X"F32D", X"0F30", X"0E15", X"F1B9", X"F2C3", X"F3B9", 
		X"0E7D", X"0D70", X"F259", X"F357", X"0EEB", X"0DD5", 
		X"F1EE", X"F2F3", X"0752", X"0E3F", X"FB6F", X"F29C", 
		X"F396", X"0EA8", X"0D97", X"F240", X"F340", X"0F12", 
		X"0DFA", X"F1E0", X"F2E7", X"F3DB", X"0E5E", X"0D52", 
		X"F28A", X"F385", X"0EB6", X"0DA4", X"F230", X"F331", 
		X"0F13", X"0DFA", X"F1D4", X"F2DC", X"F3D0", X"0E54", 
		X"0D49", X"F286", X"F381", X"0EA2", X"0D92", X"F241", 
		X"F341", X"0EFF", X"0DE8", X"F1F6", X"F2FB", X"F5F2", 
		X"0E3D", X"0942", X"F2B1", X"F3A9", X"0E84", X"0D76", 
		X"F269", X"F366", X"0ECE", X"0DBB", X"F220", X"F322", 
		X"0BEE", X"0E02", X"F372", X"F2DE", X"F3D2", X"0E4B", 
		X"0D41", X"F299", X"F392", X"0E88", X"0D79", X"F257", 
		X"F355", X"0EC8", X"0DB5", X"F215", X"F318", X"09CF", 
		X"0DF3", X"F54E", X"F2DB", X"F3D0", X"0E26", X"0D1E", 
		X"F2B1", X"F3A8", X"0E65", X"0D59", X"F280", X"F37B", 
		X"0EA2", X"0D92", X"F24D", X"F34C", X"0ED0", X"0DBD", 
		X"F21B", X"F31E", X"0707", X"0DEA", X"F563", X"F2F0", 
		X"F3E3", X"0E18", X"0D12", X"F2C3", X"F3BA", X"0E48", 
		X"0D3E", X"F2A5", X"F39D", X"0E74", X"0D67", X"F282", 
		X"F37D", X"0E9E", X"0D8E", X"F25E", X"F35C", X"0EC8", 
		X"0DB5", X"F239", X"F339", X"09B5", X"0DCF", X"F217", 
		X"F31A", X"F5FF", X"0DEB", X"FBAD", X"F2FC", X"F3EE", 
		X"0E08", X"0D03", X"F2DF", X"F3D3", X"0E26", X"0D1F", 
		X"F2C2", X"F3B8", X"0E37", X"0D2E", X"F2B7", X"F3AE", 
		X"0E54", X"0D49", X"F2A7", X"F3A0", X"0E6E", X"0D62", 
		X"F295", X"F38F", X"0E86", X"0D78", X"F281", X"F37C", 
		X"0E90", X"0D81", X"F271", X"F36D", X"0E9C", X"0D8C", 
		X"F262", X"F35F", X"0D36", X"0D98", X"F254", X"F352", 
		X"0B88", X"0D98", X"F259", X"F357", X"0992", X"0DA3", 
		X"F259", X"F357", X"06E8", X"0DAB", X"F257", X"F355", 
		X"FE21", X"0DB2", X"F254", X"F352", X"FDF0", X"0DAB", 
		X"F253", X"F352", X"FDD8", X"0DA5", X"F255", X"F353", 
		X"FDCD", X"0DA1", X"F257", X"F355", X"FDC8", X"0D9D", 
		X"F269", X"F366", X"06D8", X"0D96", X"F278", X"F374", 
		X"0985", X"0D8C", X"F285", X"F380", X"0B7B", X"0D82", 
		X"F291", X"F38B", X"0D17", X"0D77", X"F29D", X"F396", 
		X"0E6B", X"0D5F", X"F2AC", X"F3A4", X"0E54", X"0D49", 
		X"F2BD", X"F3B4", X"0E3E", X"0D35", X"F2D0", X"F3C5", 
		X"0E1B", X"0D15", X"F2E6", X"F3DA", X"0DFB", X"0CF7", 
		X"F2FE", X"F3F0", X"0DDD", X"0CDB", X"F317", X"F408", 
		X"0DC0", X"0CC0", X"F331", X"F41F", X"0D96", X"FBEE", 
		X"F35D", X"F629", X"0D79", X"F288", X"F383", X"0952", 
		X"0D58", X"F2AF", X"F3A7", X"0E40", X"0D37", X"F2D3", 
		X"F3C9", X"0E1B", X"0D15", X"F2F7", X"F3EA", X"0DE9", 
		X"0CE6", X"F31D", X"F40D", X"0DBA", X"0CBA", X"F345", 
		X"F432", X"0D8C", X"05EE", X"F36D", X"F635", X"0D5F", 
		X"F2AB", X"F3A3", X"0CCD", X"0D30", X"F2E2", X"F3D6", 
		X"0E04", X"0D00", X"F316", X"F406", X"0DD0", X"0CCF", 
		X"F348", X"F435", X"0D9C", X"0AF8", X"F379", X"F462", 
		X"0D5B", X"F2B6", X"F3AD", X"0CBA", X"0D1D", X"F2EE", 
		X"F3E2", X"0DE4", X"0CE2", X"F327", X"F416", X"0DA6", 
		X"0CA8", X"F35F", X"F44A", X"0D5C", X"F608", X"F3A8", 
		X"0923", X"0D1F", X"F2F9", X"F3EB", X"0DE3", X"0CE1", 
		X"F33D", X"F42B", X"0D9F", X"0CA2", X"F37F", X"F467", 
		X"0D4F", X"F453", X"F3C2", X"0CA0", X"0D02", X"F314", 
		X"F405", X"0DB7", X"0CB8", X"F35C", X"F447", X"0D6A", 
		X"08CC", X"F3A2", X"F8C3", X"0D1E", X"F303", X"F3F5", 
		X"0DD2", X"0CD1", X"F357", X"F443", X"0D7F", X"0C84", 
		X"F3A7", X"F48D", X"0D2C", X"F303", X"F3F5", X"0DDD", 
		X"0CDB", X"F354", X"F440", X"0D7A", X"0C80", X"F3A6", 
		X"F48C", X"0D1C", X"F307", X"F3F8", X"0DC2", X"0CC2", 
		X"F35E", X"F449", X"0D64", X"0C6B", X"F3B3", X"F669", 
		X"0D09", X"F324", X"F414", X"0DAB", X"0CAC", X"F387", 
		X"F46F", X"0D48", X"FCA2", X"F3E4", X"08FF", X"0CE7", 
		X"F353", X"F43F", X"0D84", X"0C89", X"F3B1", X"F496", 
		X"0D14", X"F320", X"F40F", X"0DA8", X"0CAA", X"F384", 
		X"F46C", X"0D3A", X"05F8", X"F3E6", X"08E5", X"0CD0", 
		X"F35B", X"F446", X"0D62", X"0C69", X"F3BF", X"F4A3", 
		X"0CEB", X"F336", X"F424", X"0D74", X"0C7A", X"F3A0", 
		X"F487", X"0CFF", X"F497", X"F409", X"0D8B", X"0C8F", 
		X"F386", X"F46F", X"0D17", X"FC7C", X"F3FE", X"0C41", 
		X"0CA4", X"F387", X"F46F", X"0D27", X"08AC", X"F3FA", 
		X"08CB", X"0CB0", X"F381", X"F469", X"0D33", X"0C3D", 
		X"F3F3", X"FD31", X"0CBB", X"F378", X"F462", X"0D30", 
		X"0C3B", X"F3EE", X"FD00", X"0CAD", X"F378", X"F461", 
		X"0D25", X"0C31", X"F3F1", X"FCF2", X"0CA5", X"F37C", 
		X"F465", X"0D1E", X"0C2A", X"F403", X"0613", X"0C9B", 
		X"F39B", X"F482", X"0D0E", X"08A0", X"F41C", X"0A96", 
		X"0C89", X"F3B3", X"F498", X"0CFA", X"FCC7", X"F432", 
		X"0D6F", X"0C75", X"F3C8", X"F4AC", X"0CD8", X"F4D8", 
		X"F449", X"0D41", X"0C4A", X"F3E5", X"F4C7", X"0CAF", 
		X"F37F", X"F468", X"0D18", X"0C24", X"F406", X"F8E5", 
		X"0C89", X"F3B0", X"F495", X"0CEE", X"05EB", X"F440", 
		X"0D54", X"0C5C", X"F3E7", X"F4C9", X"0CBD", X"F38B", 
		X"F473", X"0D20", X"0C2C", X"F41B", X"F6B6", X"0C8A", 
		X"F3BF", X"F4A3", X"0CDF", X"05E5", X"F44F", X"0D37", 
		X"0C41", X"F3F9", X"F4D9", X"0C97", X"F3A3", X"F489", 
		X"0CEF", X"0BFF", X"F437", X"087D", X"0C53", X"F3E2", 
		X"F4C4", X"0C9E", X"F39D", X"F484", X"0CF6", X"0C05", 
		X"F43F", X"05ED", X"0C56", X"F3F6", X"F4D6", X"0CA8", 
		X"F3A9", X"F48F", X"0CFC", X"0C0A", X"F446", X"FD28", 
		X"0C59", X"F3FA", X"F4DA", X"0C9D", X"F3B0", X"F495", 
		X"0CE4", X"0BF4", X"F450", X"086B", X"0C39", X"F40A", 
		X"F4E9", X"0C7F", X"F3C3", X"F4A7", X"0CC8", X"0BDA", 
		X"F464", X"0D06", X"0C13", X"F430", X"F50C", X"0C59", 
		X"F3F8", X"F4D8", X"0C9D", X"F6E9", X"F4A0", X"0CE2", 
		X"0BF2", X"F466", X"05E0", X"0C32", X"F42B", X"F507", 
		X"0C72", X"F3ED", X"F4CE", X"0CA8", X"05E0", X"F496", 
		X"0CDF", X"0BF0", X"F45F", X"FCF4", X"0C26", X"F428", 
		X"F505", X"0C5D", X"F3F1", X"F4D1", X"0C96", X"05CF", 
		X"F49D", X"0CC3", X"0BD5", X"F478", X"084A", X"0C0B", 
		X"F44F", X"F529", X"0C3F", X"F423", X"F500", X"0C72", 
		X"F3F6", X"F4D6", X"0CA5", X"0A3E", X"F4AA", X"0CD9", 
		X"0BEA", X"F47D", X"FD0D", X"0C0E", X"F452", X"F52C", 
		X"0C34", X"F428", X"F505", X"0C5C", X"F3FF", X"F4DE", 
		X"0C86", X"0853", X"F4B7", X"0CB0", X"0BC3", X"F491", 
		X"0831", X"0BEB", X"F469", X"F541", X"0C07", X"F445", 
		X"F51F", X"0C26", X"F421", X"F4FF", X"0C46", X"F568", 
		X"F4DE", X"0C67", X"0836", X"F4BE", X"0C89", X"0BA0", 
		X"F49F", X"0B5E", X"0BC0", X"F47E", X"FC96", X"0BD5", 
		X"F46E", X"F546", X"0BF4", X"F45A", X"F533", X"0C12", 
		X"F444", X"F51F", X"0C2F", X"F42C", X"F509", X"0C4B", 
		X"F95B", X"F4F2", X"0C66", X"0A0A", X"F4DA", X"0C82", 
		X"0B99", X"F4C3", X"0C91", X"0BA7", X"F4AD", X"0802", 
		X"0BB6", X"F499", X"F925", X"0BC7", X"F486", X"F55B", 
		X"0BD9", X"F473", X"F54A", X"0BEB", X"F460", X"F539", 
		X"0BFD", X"F45B", X"F534", X"0C0D", X"F453", X"F52D", 
		X"0C1B", X"F44A", X"F524", X"0C28", X"F751", X"F51B", 
		X"0C35", X"FD7C", X"F511", X"0C41", X"082C", X"F507", 
		X"0C4D", X"0B68", X"F4FD", X"0C4D", X"0B68", X"F4F5", 
		X"0C4E", X"0B69", X"F4EF", X"0C51", X"0B6B", X"F4EA", 
		X"0C54", X"0B6F", X"F4E5", X"0C58", X"0B72", X"F4E0", 
		X"0B16", X"0B76", X"F4DC", X"09A0", X"0B7A", X"F4E5", 
		X"09A4", X"0B7B", X"F4EB", X"09A5", X"0B7A", X"F4F0", 
		X"09A5", X"0B79", X"F4F4", X"09A4", X"0B77", X"F4F8", 
		X"09A2", X"0B75", X"F4FB", X"09A0", X"0B72", X"F4FE", 
		X"099E", X"0B70", X"F501", X"0B04", X"0B61", X"F506", 
		X"0C39", X"0B55", X"F50D", X"0C2C", X"0B4A", X"F515", 
		X"0C21", X"0B3F", X"F51E", X"0C16", X"0B35", X"F527", 
		X"0C0B", X"0B2B", X"F52F", X"0BF5", X"059C", X"F547", 
		X"0BE9", X"F9A9", X"F55C", X"0BDC", X"F5F8", X"F56F", 
		X"0BCD", X"F4AD", X"F580", X"0BBD", X"F4BF", X"F590", 
		X"0BAD", X"F4D0", X"F5A0", X"0B9C", X"F4E0", X"F5B0", 
		X"0B80", X"F4F4", X"F5C1", X"0B66", X"F508", X"FCCA", 
		X"0B4D", X"F51D", X"0966", X"0B34", X"F533", X"0BFC", 
		X"0B1D", X"F548", X"0BE3", X"09A1", X"F55E", X"0BCA", 
		X"FD9C", X"F574", X"0BB2", X"F4C4", X"F595", X"0B97", 
		X"F4E6", X"F5B5", X"0B7B", X"F506", X"F5D2", X"0B5E", 
		X"F524", X"F97E", X"0B41", X"F542", X"095C", X"0B23", 
		X"F55F", X"0BE3", X"0B06", X"F57C", X"0BC4", X"FE15", 
		X"F598", X"0B99", X"F4E7", X"F5B6", X"0B71", X"F509", 
		X"F5D5", X"0B4A", X"F52B", X"F976", X"0B24", X"F54D", 
		X"0AA2", X"0AFF", X"F570", X"0BB5", X"07D4", X"F592", 
		X"0B8F", X"F639", X"F5B4", X"0B5D", X"F50B", X"F5D7", 
		X"0B2E", X"F533", X"FC9C", X"0B01", X"F55B", X"0BB0", 
		X"0AD6", X"F583", X"0B82", X"F9CD", X"F5AB", X"0B55", 
		X"F505", X"F5D2", X"0B29", X"F52F", X"F779", X"0AFE", 
		X"F559", X"0BA1", X"0AC8", X"F590", X"0B73", X"F7D9", 
		X"F5C4", X"0B44", X"F52A", X"F5F4", X"0B14", X"F55D", 
		X"04F8", X"0AE4", X"F58D", X"0B8C", X"07BB", X"F5BD", 
		X"0B59", X"F520", X"F5EB", X"0B27", X"F551", X"F797", 
		X"0AEA", X"F583", X"0B87", X"0AB1", X"F5B6", X"0B4B", 
		X"F51D", X"F5E8", X"0B11", X"F553", X"F796", X"0AD9", 
		X"F589", X"0B77", X"0AA2", X"F5BD", X"0B3D", X"F526", 
		X"F5F1", X"0B04", X"F569", X"F98E", X"0ACA", X"F5A9", 
		X"0B64", X"0572", X"F5E5", X"0B25", X"F559", X"F620", 
		X"0AE8", X"F596", X"08EF", X"0AAB", X"F5D1", X"0B41", 
		X"F68F", X"F60B", X"0B02", X"F580", X"F7BD", X"0AC4", 
		X"F5BB", X"0B4F", X"0568", X"F5F8", X"0B06", X"F56F", 
		X"F634", X"0ABF", X"F5AF", X"0B4E", X"092A", X"F5EE", 
		X"0B07", X"F567", X"F62D", X"0AC1", X"F5A9", X"0A22", 
		X"0A7E", X"F5E9", X"0B0A", X"F562", X"F628", X"0ABA", 
		X"F5B2", X"0A1B", X"0A77", X"F5FD", X"0B00", X"F581", 
		X"F645", X"0AB7", X"F5CB", X"0B41", X"0924", X"F612", 
		X"0AF5", X"F594", X"F656", X"0AAB", X"F5DC", X"0B33", 
		X"0789", X"F621", X"0AE7", X"F5A4", X"F665", X"0A92", 
		X"F5ED", X"0B0F", X"FA3C", X"F635", X"0ABB", X"F5BD", 
		X"04A8", X"0A6B", X"F608", X"0AE8", X"F58F", X"F652", 
		X"0A97", X"F5DC", X"0B17", X"08FF", X"F627", X"0AC4", 
		X"F5AF", X"F670", X"0A74", X"F608", X"0AF0", X"F6DC", 
		X"F65B", X"0A9B", X"F5EF", X"09F0", X"0903", X"F641", 
		X"0ABF", X"F5D2", X"F7FD", X"0A6A", X"F624", X"0AE2", 
		X"F5B3", X"F673", X"0A8B", X"F606", X"0B04", X"076E", 
		X"F656", X"0AAC", X"F5E7", X"FCDA", X"0A4C", X"F63A", 
		X"0AB9", X"F5CE", X"F68C", X"0A5B", X"F624", X"0ACA", 
		X"F6F6", X"F678", X"0A6D", X"F610", X"0ADD", X"0538", 
		X"F665", X"0A7F", X"F5FC", X"06D5", X"0A25", X"F652", 
		X"0A93", X"F5F5", X"F9E0", X"0A35", X"F655", X"0AA0", 
		X"F5F4", X"F6B0", X"0A41", X"F652", X"0AAA", X"F5F0", 
		X"F6AC", X"0A49", X"F64D", X"0AB3", X"F5EB", X"F6A7", 
		X"0A51", X"F648", X"0ABA", X"F89E", X"F6A1", X"0A58", 
		X"F642", X"0AB7", X"FA8D", X"F69D", X"0A4B", X"F641", 
		X"0AAC", X"FA87", X"F69E", X"0A43", X"F643", X"0AA4", 
		X"FA86", X"F6A2", X"0A3C", X"F648", X"0A9D", X"FA87", 
		X"F6A6", X"0A35", X"F64C", X"0A97", X"FA8A", X"F6AB", 
		X"0A2F", X"F652", X"0A86", X"F8A0", X"F6B2", X"0A16", 
		X"F65C", X"0A6E", X"F604", X"F6BE", X"0A01", X"F66A", 
		X"0A5A", X"F614", X"F6CD", X"09EE", X"F67A", X"0A47", 
		X"F625", X"F9E7", X"09DC", X"F68A", X"0A34", X"F636", 
		X"0436", X"09CA", X"F6A6", X"0A20", X"F65C", X"0A77", 
		X"FE71", X"F6C7", X"0A06", X"F67C", X"0A5B", X"F62E", 
		X"F6E5", X"09EA", X"F69A", X"0A3D", X"F64C", X"FA0D", 
		X"09CD", X"F6B7", X"0A1F", X"F66A", X"0815", X"070B", 
		X"F6D3", X"0A01", X"F687", X"0A4A", X"F76A", X"F6F0", 
		X"09D1", X"F6A8", X"0A1A", X"F65E", X"042A", X"09A5", 
		X"F6CC", X"09EE", X"F685", X"0A3A", X"F8D1", X"F6F1", 
		X"09C4", X"F6AB", X"0A0F", X"F663", X"FCAC", X"099B", 
		X"F6D2", X"09E4", X"F68B", X"0A30", X"F8E2", X"F703", 
		X"09B9", X"F6C7", X"0A00", X"F688", X"0666", X"06F0", 
		X"F6FC", X"09CE", X"F6BD", X"0A14", X"F67D", X"F87D", 
		X"099A", X"F6F0", X"09DF", X"F6B1", X"0A25", X"F902", 
		X"F722", X"09AA", X"F6E3", X"09EE", X"F6A3", X"07DA", 
		X"04F3", X"F716", X"09A7", X"F6DA", X"09E3", X"F69D", 
		X"0645", X"06D0", X"F713", X"09A0", X"F6D9", X"09DD", 
		X"F69D", X"0405", X"0836", X"F714", X"099C", X"F6DA", 
		X"09DA", X"F69F", X"FCBD", X"095C", X"F716", X"0999", 
		X"F6DD", X"09CC", X"F6AF", X"03FF", X"06C4", X"F72F", 
		X"0989", X"F6FF", X"09C3", X"F6CC", X"07B8", X"FF08", 
		X"F748", X"097A", X"F716", X"09B2", X"F6E3", X"09EB", 
		X"F934", X"F75C", X"0968", X"F72A", X"099F", X"F6F7", 
		X"09D7", X"F6C3", X"F76F", X"0954", X"F748", X"097F", 
		X"F715", X"09AD", X"F6E3", X"079C", X"FEDE", X"F75F", 
		X"0952", X"F731", X"0981", X"F702", X"09B1", X"F6D2", 
		X"FA51", X"092B", X"F751", X"095A", X"F723", X"098A", 
		X"F6F5", X"08B3", X"FB02", X"F772", X"0935", X"F746", 
		X"095B", X"F724", X"098B", X"F700", X"0780", X"FB1C", 
		X"F785", X"0930", X"F761", X"095C", X"F73B", X"0988", 
		X"F713", X"0780", X"FB2E", X"F795", X"0929", X"F76F", 
		X"0953", X"F748", X"097E", X"F720", X"0778", X"FB37", 
		X"F7A1", X"091E", X"F77A", X"093E", X"F755", X"0960", 
		X"F730", X"0983", X"F70C", X"FA76", X"07DA", X"F791", 
		X"0916", X"F76F", X"0939", X"F74C", X"095D", X"F72A", 
		X"0753", X"FB2D", X"F7AE", X"08F3", X"F78D", X"0916", 
		X"F76B", X"093A", X"F749", X"095E", X"F727", X"03B4", 
		X"FEF4", X"F7B7", X"08EB", X"F7A0", X"090C", X"F787", 
		X"092D", X"F76D", X"094D", X"F752", X"0748", X"F99D", 
		X"F7DA", X"08DB", X"F7C0", X"08F9", X"F7A5", X"0917", 
		X"F789", X"0936", X"F76D", X"0955", X"F751", X"FAAC", 
		X"066D", X"F7D9", X"08E1", X"F7BD", X"08F5", X"F7A3", 
		X"090B", X"F78A", X"0922", X"F772", X"0939", X"F759", 
		X"FCFF", X"0497", X"F7E4", X"08BA", X"F7CE", X"08D1", 
		X"F7B7", X"08E9", X"F7A0", X"0901", X"F789", X"0919", 
		X"F772", X"05AC", X"FB61", X"F7FC", X"089D", X"F7E7", 
		X"08B4", X"F7D1", X"08C3", X"F7BC", X"08D2", X"F7A8", 
		X"08E3", X"F795", X"08F4", X"F782", X"080D", X"F87A", 
		X"FCD9", X"0466", X"F7FE", X"087F", X"F7ED", X"0891", 
		X"F7DC", X"08A3", X"F7CA", X"08B5", X"F7B9", X"08C7", 
		X"F7A8", X"08D9", X"F796", X"07F5", X"F88C", X"035A", 
		X"FB63", X"F93E", X"0616", X"F816", X"086E", X"F80D", 
		X"087D", X"F803", X"088B", X"F7F9", X"0899", X"F7EE", 
		X"08A6", X"F7E3", X"08B4", X"F7D7", X"08C1", X"F7CC", 
		X"08CE", X"F7C0", X"06D1", X"F8BA", X"FD15", X"FF8D", 
		X"F844", X"074B", X"F839", X"085A", X"F82D", X"085E", 
		X"F823", X"0863", X"F81A", X"0868", X"F812", X"086E", 
		X"F80A", X"0874", X"F802", X"087B", X"F7FA", X"0882", 
		X"F7F3", X"0889", X"F7EC", X"0890", X"F7E5", X"0897", 
		X"F7DE", X"07B0", X"F7D6", X"0546", X"FA00", X"FCF6", 
		X"FED6", X"F978", X"05DD", X"F85C", X"05DD", X"F85F", 
		X"0718", X"F862", X"081B", X"F863", X"0820", X"F863", 
		X"0823", X"F862", X"0826", X"F862", X"0829", X"F861", 
		X"082C", X"F85F", X"082E", X"F85E", X"0831", X"F85C", 
		X"0833", X"F85B", X"0835", X"F859", X"0837", X"F857", 
		X"0839", X"F856", X"083B", X"F854", X"0834", X"F854", 
		X"082F", X"F854", X"082A", X"F855", X"0825", X"F857", 
		X"0821", X"F859", X"081E", X"F85B", X"081A", X"F85E", 
		X"0817", X"F860", X"0813", X"F863", X"0810", X"F866", 
		X"080D", X"F868", X"080A", X"F86B", X"0807", X"F86E", 
		X"0803", X"F871", X"0800", X"F87D", X"07FC", X"F887", 
		X"07F6", X"F891", X"07F0", X"F89A", X"07EA", X"F8A3", 
		X"07E3", X"F8AB", X"07DB", X"F8B3", X"07D4", X"F8BA", 
		X"07CD", X"F8C2", X"07C5", X"F8C9", X"07BE", X"F8D1", 
		X"07B6", X"F8D8", X"06C1", X"F8DF", X"059E", X"F8E7", 
		X"041E", X"F9F5", X"00DF", X"FD48", X"FA81", X"04F1", 
		X"F879", X"0725", X"F884", X"07F3", X"F88F", X"07E6", 
		X"F89A", X"07D8", X"F8A5", X"07CB", X"F8B0", X"07BE", 
		X"F8BC", X"07B1", X"F8C7", X"07A5", X"F8D3", X"0798", 
		X"F8DE", X"078C", X"F8EA", X"077F", X"F8F5", X"0773", 
		X"F901", X"0567", X"FA0A", X"FF57", X"02EB", X"F8A2", 
		X"06F6", X"F8B6", X"07BF", X"F8C9", X"07B0", X"F8DC", 
		X"07A0", X"F8ED", X"0791", X"F8FE", X"0781", X"F90E", 
		X"0770", X"F91F", X"0760", X"F92E", X"03F9", X"FB79", 
		X"FAC5", X"04C7", X"F8D6", X"07B0", X"F8E6", X"079F", 
		X"F8F7", X"078E", X"F906", X"077D", X"F916", X"076C", 
		X"F926", X"0753", X"F936", X"073C", X"F948", X"00A8", 
		X"02E8", X"F8E6", X"0789", X"F8F9", X"0772", X"F90D", 
		X"075D", X"F920", X"0747", X"F934", X"0732", X"F947", 
		X"071D", X"F95A", X"0020", X"02D4", X"F8FC", X"076C", 
		X"F910", X"0756", X"F924", X"0741", X"F938", X"072C", 
		X"F94B", X"0717", X"F95E", X"051C", X"FB95", X"F9EF", 
		X"0691", X"F92D", X"0745", X"F947", X"072D", X"F960", 
		X"0715", X"F978", X"06FD", X"F990", X"FC74", X"0485", 
		X"F93F", X"073F", X"F956", X"0726", X"F96E", X"070D", 
		X"F985", X"06F4", X"F99C", X"03C2", X"FD9C", X"F94B", 
		X"0734", X"F962", X"071A", X"F979", X"0701", X"F990", 
		X"06E2", X"F9A8", X"03AD", X"02C0", X"F95B", X"070E", 
		X"F975", X"06F0", X"F990", X"06D3", X"F9A9", X"05E7", 
		X"FBC7", X"FA33", X"0703", X"F97B", X"06E5", X"F996", 
		X"06C9", X"F9B0", X"06AD", X"F9CA", X"FC86", X"0557", 
		X"F983", X"06DC", X"F99E", X"06C0", X"F9B8", X"06A4", 
		X"F9D2", X"0383", X"0431", X"F98C", X"06C5", X"F9A9", 
		X"06A3", X"F9C5", X"0683", X"FABD", X"FB44", X"06C3", 
		X"F9A2", X"06A3", X"F9C0", X"0683", X"F9DD", X"04A7", 
		X"0269", X"F99F", X"06A4", X"F9BD", X"0684", X"F9DB", 
		X"0665", X"F9F8", X"FC91", X"05EA", X"F9BB", X"0686", 
		X"F9D9", X"0666", X"F9F6", X"0582", X"FD7A", X"F9B9", 
		X"0680", X"F9DF", X"0661", X"FA04", X"057E", X"FD92", 
		X"F9D3", X"067C", X"F9F6", X"065A", X"FA17", X"0578", 
		X"FDA5", X"F9E5", X"0671", X"FA06", X"064E", X"FA27", 
		X"056E", X"FDAF", X"F9F4", X"0663", X"FA15", X"0640", 
		X"FA35", X"0562", X"FDB6", X"FA02", X"0654", X"FA23", 
		X"0632", X"FA43", X"0556", X"FDBC", X"FA10", X"063F", 
		X"FA32", X"0617", X"FA53", X"0034", X"0593", X"FA26", 
		X"061B", X"FA48", X"05F6", X"FC2C", X"FA1C", X"0621", 
		X"FA40", X"05FC", X"FA62", X"0319", X"04B0", X"FA38", 
		X"0603", X"FA5B", X"05DE", X"FB42", X"FAE8", X"0609", 
		X"FA54", X"05E5", X"FA77", X"0432", X"03A3", X"FA4E", 
		X"05EB", X"FA71", X"05C7", X"FB53", X"FA4F", X"05EB", 
		X"FA78", X"05C6", X"FAA0", X"FBE7", X"05ED", X"FA82", 
		X"05C6", X"FAA8", X"00BB", X"0546", X"FA88", X"05C4", 
		X"FAAD", X"0421", X"0397", X"FA8E", X"05C0", X"FAB3", 
		X"0599", X"FDEA", X"FA93", X"05BB", X"FAB7", X"0594", 
		X"FB97", X"FA98", X"05B6", X"FABC", X"0590", X"FAE0", 
		X"FC1B", X"05B1", X"FAC1", X"0585", X"FAE6", X"FC1D", 
		X"059B", X"FACA", X"0571", X"FAF0", X"FB58", X"0589", 
		X"FAD6", X"0560", X"FBAF", X"FABD", X"0578", X"FAE4", 
		X"0550", X"FC98", X"FACC", X"0568", X"FAF2", X"0540", 
		X"FDE8", X"FADB", X"0558", X"FB01", X"0530", X"01ED", 
		X"FAEA", X"0548", X"FB10", X"0481", X"0339", X"FAF9", 
		X"0538", X"FB1F", X"03B4", X"04B4", X"FB0F", X"0522", 
		X"FB3A", X"FBA3", X"0537", X"FB2E", X"050E", X"FE15", 
		X"FB20", X"0521", X"FB48", X"02B7", X"04A2", X"FB3A", 
		X"0508", X"FB61", X"FBC7", X"0519", X"FB53", X"04EF", 
		X"FE2C", X"FB44", X"04FF", X"FB6B", X"02A7", X"0483", 
		X"FB5D", X"04E6", X"FB83", X"FBE6", X"04F5", X"FB75", 
		X"04CC", X"FE3A", X"FB67", X"04DB", X"FB8D", X"00B8", 
		X"04E0", X"FB81", X"04B3", X"FE2E", X"FB77", X"04BA", 
		X"FB9F", X"FD99", X"04C1", X"FB96", X"0497", X"01B3", 
		X"FB8E", X"049E", X"FBB6", X"FCC0", X"04A6", X"FBAE", 
		X"047C", X"02CE", X"FBA7", X"0483", X"FBCE", X"FC2B", 
		X"048A", X"FBC8", X"03D9", X"037A", X"FBC1", X"0467", 
		X"FBE8", X"FBBB", X"046E", X"FBE2", X"0321", X"03F7", 
		X"FBE1", X"044B", X"FE59", X"FBE3", X"044F", X"FC0C", 
		X"FBE5", X"0451", X"FC0E", X"00BC", X"0452", X"FC0E", 
		X"0428", X"02A1", X"FC0F", X"0428", X"FCC0", X"FC0F", 
		X"0428", X"FC36", X"FD2B", X"0428", X"FC37", X"02F4", 
		X"03B4", X"FC38", X"03FE", X"FE8A", X"FC39", X"03FD", 
		X"FC5F", X"FC3A", X"03FC", X"FC60", X"00B9", X"03FA", 
		X"FC61", X"03D2", X"026B", X"FC63", X"03CC", X"FE92", 
		X"FC67", X"03C3", X"FD09", X"FC6B", X"03BA", X"FC92", 
		X"FC71", X"03B2", X"FC98", X"FD71", X"03AA", X"FC9E", 
		X"006E", X"03A2", X"FCA5", X"028E", X"039A", X"FCAD", 
		X"0372", X"02B7", X"FCB5", X"0369", X"0140", X"FCBD", 
		X"0361", X"FDDC", X"FCC5", X"0358", X"FCEA", X"FCCE", 
		X"034F", X"FCF3", X"FD3C", X"0345", X"FCFC", X"FE5D", 
		X"0338", X"FD09", X"FDCB", X"032D", X"FD19", X"FDD8", 
		X"0320", X"FD28", X"FDE5", X"0312", X"FD37", X"FDF0", 
		X"0304", X"FD46", X"FDFC", X"02F4", X"FD55", X"FE07", 
		X"02E5", X"FD64", X"FE12", X"02D4", X"FD73", X"FE1E", 
		X"02C3", X"FD83", X"FE2A", X"02B2", X"FD93", X"FE36", 
		X"02A0", X"FDA3", X"FE42", X"028E", X"FDB4", X"FE4F", 
		X"027A", X"FDC6", X"FE5C", X"0266", X"FDD8", X"FE12", 
		X"024D", X"FDEC", X"FDE0", X"0234", X"FE49", X"FDF6", 
		X"021A", X"FF32", X"FE0E", X"0200", X"0139", X"FE27", 
		X"01E5", X"01B7", X"FE42", X"0150", X"01CF", X"FE5E", 
		X"003D", X"01AF", X"FE7C", X"FEE5", X"018D", X"FE9C", 
		X"FE9B", X"0168", X"FEC0", X"FEC1", X"013E", X"FF40", 
		X"FEED", X"010E", X"005C", X"FF22", X"00D2", X"0092", 
		X"FF6C", X"0066", X"002C");

	constant sound2 : sound2_type :=	 (
		X"0000", X"0CA1", X"11BA", X"1555", X"181B", X"1A4C", 
		X"1C00", X"1D4A", X"1E30", X"1EBA", X"1EE7", X"1EBB", 
		X"1E32", X"1D4D", X"1C02", X"1A4F", X"181A", X"1555", 
		X"11B1", X"0C9B", X"FAD8", X"F1FF", X"ED54", X"E9EF", 
		X"E759", X"E547", X"E3B7", X"E28B", X"E1C7", X"E15F", 
		X"E155", X"E1A8", X"E257", X"E36E", X"E4E6", X"E6DF", 
		X"E967", X"EC8F", X"F0F1", X"F806", X"0B0F", X"10B0", 
		X"1481", X"1767", X"19AE", X"1B73", X"1CCA", X"1DBA", 
		X"1E4B", X"1E7F", X"1E56", X"1DD0", X"1CEB", X"1B9F", 
		X"19E8", X"17AC", X"14DB", X"1121", X"0BCF", X"F92D", 
		X"F17C", X"ED08", X"E9D0", X"E746", X"E554", X"E3D0", 
		X"E2BA", X"E20C", X"E1BC", X"E1CB", X"E23A", X"E307", 
		X"E440", X"E5DF", X"E809", X"EABB", X"EE58", X"F350", 
		X"04D0", X"0DCC", X"1263", X"15B7", X"184B", X"1A4F", 
		X"1BD8", X"1CF8", X"1DB2", X"1E0D", X"1E09", X"1DA7", 
		X"1CE6", X"1BBD", X"1A2C", X"181A", X"157C", X"120A", 
		X"0D50", X"01FB", X"F2FA", X"EE19", X"EAAF", X"E803", 
		X"E5F9", X"E463", X"E33D", X"E282", X"E227", X"E22E", 
		X"E296", X"E35E", X"E494", X"E631", X"E85B", X"EB10", 
		X"EEB6", X"F3C9", X"05E0", X"0E0E", X"1281", X"15BF", 
		X"1841", X"1A33", X"1BAD", X"1CBA", X"1D64", X"1DAB", 
		X"1D93", X"1D1B", X"1C3F", X"1AF9", X"1945", X"1708", 
		X"142F", X"1060", X"0AC6", X"F7D0", X"F107", X"ECD4", 
		X"E9C7", X"E760", X"E58F", X"E42D", X"E33D", X"E2B0", 
		X"E287", X"E2C1", X"E35B", X"E462", X"E5CF", X"E7C2", 
		X"EA37", X"ED7F", X"F1DF", X"FA2B", X"0BEE", X"110A", 
		X"1495", X"1749", X"1960", X"1AF9", X"1C20", X"1CE0", 
		X"1D3C", X"1D37", X"1CD0", X"1C03", X"1AD0", X"1927", 
		X"16F9", X"1431", X"1077", X"0B0B", X"F85E", X"F15C", 
		X"ED21", X"EA11", X"E7AB", X"E5DD", X"E480", X"E396", 
		X"E310", X"E2F1", X"E336", X"E3DD", X"E4F4", X"E674", 
		X"E880", X"EB15", X"EE92", X"F35F", X"040D", X"0D5B", 
		X"11E7", X"152A", X"17AC", X"1998", X"1B0A", X"1C0C", 
		X"1CA7", X"1CDD", X"1CB0", X"1C20", X"1B25", X"19C0", 
		X"17DA", X"156B", X"1233", X"0DD3", X"0588", X"F418", 
		X"EF05", X"EB8F", X"E8E3", X"E6DF", X"E555", X"E444", 
		X"E39A", X"E359", X"E37E", X"E407", X"E4FF", X"E65F", 
		X"E849", X"EAB7", X"EDFD", X"F266", X"FB51", X"0C29", 
		X"110C", X"1476", X"170F", X"190C", X"1A8B", X"1B96", 
		X"1C39", X"1C74", X"1C4B", X"1BBD", X"1AC3", X"195D", 
		X"1774", X"14FD", X"11B7", X"0D37", X"039F", X"F39B", 
		X"EED8", X"EB71", X"E8E9", X"E6F1", X"E582", X"E47F", 
		X"E3ED", X"E3C1", X"E3FC", X"E4A2", X"E5B0", X"E73C", 
		X"E940", X"EBF5", X"EF75", X"F4BB", X"0694", X"0DFD", 
		X"1230", X"1541", X"1797", X"195E", X"1AA9", X"1B86", 
		X"1BF8", X"1C04", X"1BAA", X"1AE5", X"19B4", X"1808", 
		X"15D7", X"12EF", X"0F12", X"08D9", X"F65F", X"F085", 
		X"ECCA", X"E9F8", X"E7DC", X"E647", X"E523", X"E473", 
		X"E42B", X"E44D", X"E4DA", X"E5D0", X"E742", X"E92C", 
		X"EBC2", X"EF18", X"F406", X"049D", X"0D3A", X"1199", 
		X"14BD", X"171E", X"18ED", X"1A3D", X"1B1C", X"1B8F", 
		X"1B9B", X"1B3E", X"1A75", X"193F", X"1789", X"154B", 
		X"125B", X"0E4A", X"0793", X"F566", X"F01E", X"EC85", 
		X"E9E2", X"E7D8", X"E65E", X"E555", X"E4BF", X"E494", 
		X"E4D2", X"E57F", X"E698", X"E834", X"EA4E", X"ED28", 
		X"F0E9", X"F6FE", X"0944", X"0F15", X"12D2", X"1594", 
		X"17AF", X"193D", X"1A55", X"1AFC", X"1B39", X"1B0C", 
		X"1A74", X"196E", X"17EE", X"15ED", X"133F", X"0FB3", 
		X"0A4D", X"F855", X"F1C6", X"EDC6", X"EAE8", X"E8B3", 
		X"E717", X"E5F1", X"E542", X"E4FD", X"E526", X"E5BD", 
		X"E6C1", X"E847", X"EA4B", X"ED09", X"F0A2", X"F652", 
		X"0863", X"0E88", X"125A", X"1526", X"1745", X"18D7", 
		X"19EF", X"1A95", X"1ACF", X"1A9F", X"1A01", X"18F4", 
		X"176A", X"155A", X"12A2", X"0EE6", X"0926", X"F6FC", 
		X"F130", X"ED71", X"EABC", X"E8A9", X"E72A", X"E621", 
		X"E58E", X"E568", X"E5AF", X"E662", X"E791", X"E935", 
		X"EB7B", X"EE6C", X"F2A1", X"FA0B", X"0B19", X"0FF9", 
		X"1350", X"15CB", X"17A9", X"1901", X"19E2", X"1A55", 
		X"1A5A", X"19F2", X"191C", X"17CD", X"15FF", X"138E", 
		X"1055", X"0B9F", X"FB87", X"F319", X"EEE6", X"EBE8", 
		X"E9A0", X"E7F8", X"E6CA", X"E617", X"E5D2", X"E5FC", 
		X"E699", X"E7A5", X"E937", X"EB4E", X"EE15", X"F203", 
		X"F85A", X"09F5", X"0F33", X"12AB", X"153A", X"1725", 
		X"1887", X"1970", X"19E7", X"19F1", X"198C", X"18B8", 
		X"1769", X"1599", X"1324", X"0FE1", X"0B0B", X"FA57", 
		X"F2E9", X"EECE", X"EBEB", X"E9BA", X"E826", X"E70C", 
		X"E66D", X"E63D", X"E67D", X"E732", X"E859", X"E9FF", 
		X"EC4C", X"EF4C", X"F3AF", X"FD01", X"0BCD", X"103E", 
		X"1358", X"15A5", X"1758", X"188A", X"1944", X"198D", 
		X"1968", X"18D1", X"17C7", X"163C", X"1425", X"1159", 
		X"0D6C", X"06BF", X"F592", X"F0AA", X"ED51", X"EAE5", 
		X"E912", X"E7D0", X"E706", X"E6AC", X"E6C5", X"E753", 
		X"E852", X"E9D9", X"EBE6", X"EEBE", X"F294", X"F921", 
		X"0A61", X"0F42", X"128A", X"14F4", X"16BE", X"1800", 
		X"18C9", X"191F", X"1905", X"1879", X"1779", X"15F8", 
		X"13EA", X"111E", X"0D48", X"06AC", X"F5AE", X"F0D4", 
		X"ED86", X"EB25", X"E95C", X"E823", X"E761", X"E716", 
		X"E73C", X"E7D7", X"E8E6", X"EA82", X"ECA8", X"EFA6", 
		X"F3C8", X"FC4C", X"0B62", X"0FC8", X"12D5", X"1513", 
		X"16B9", X"17D8", X"1881", X"18B6", X"187A", X"17CA", 
		X"16A3", X"14F4", X"12AD", X"0F8D", X"0B10", X"FB71", 
		X"F38C", X"EF90", X"ECB3", X"EAA1", X"E91C", X"E821", 
		X"E79B", X"E789", X"E7E9", X"E8C4", X"EA18", X"EC04", 
		X"EE90", X"F210", X"F7D9", X"08E1", X"0E30", X"1196", 
		X"1411", X"15E1", X"1726", X"17F1", X"1845", X"1827", 
		X"1796", X"168B", X"1501", X"12E2", X"0FF7", X"0BDB", 
		X"0267", X"F490", X"F046", X"ED5C", X"EB37", X"E9A4", 
		X"E89E", X"E80D", X"E7F4", X"E851", X"E922", X"EA6F", 
		X"EC57", X"EEDE", X"F27B", X"F833", X"0901", X"0E25", 
		X"1175", X"13DF", X"15A0", X"16D9", X"1793", X"17D9", 
		X"17AC", X"170A", X"15EC", X"144B", X"1206", X"0EF5", 
		X"0A72", X"FA72", X"F38C", X"EFB6", X"ED0B", X"EB0F", 
		X"E9B0", X"E8D1", X"E867", X"E875", X"E8FA", X"E9F6", 
		X"EB74", X"ED98", X"F071", X"F4AE", X"01B9", X"0B7A", 
		X"0F89", X"125C", X"146D", X"15E5", X"16DC", X"1758", 
		X"175F", X"16F3", X"160F", X"14A7", X"12B0", X"0FF8", 
		X"0C2B", X"0517", X"F585", X"F127", X"EE25", X"EC01", 
		X"EA78", X"E970", X"E8E8", X"E8D6", X"E93A", X"EA1C", 
		X"EB7A", X"ED69", X"F025", X"F3EB", X"FB63", X"0A81", 
		X"0ECE", X"11BC", X"13DB", X"1560", X"165F", X"16E3", 
		X"16F2", X"168C", X"15AB", X"144C", X"1253", X"0FA7", 
		X"0BDC", X"0458", X"F57D", X"F130", X"EE52", X"EC3E", 
		X"EABD", X"E9CA", X"E94F", X"E94D", X"E9C5", X"EAB4", 
		X"EC26", X"EE3F", X"F110", X"F54C", X"037C", X"0B79", 
		X"0F52", X"11FE", X"13EF", X"154A", X"1623", X"1683", 
		X"166D", X"15DF", X"14D7", X"134A", X"1117", X"0E17", 
		X"097F", X"F9CF", X"F3B3", X"F024", X"EDAC", X"EBDD", 
		X"EAA8", X"E9F1", X"E9B2", X"E9EB", X"EAA1", X"EBD2", 
		X"ED8F", X"F00A", X"F372", X"F967", X"0923", X"0DBF", 
		X"10C2", X"12EC", X"1477", X"1578", X"15FF", X"160D", 
		X"15A6", X"14C2", X"135E", X"115D", X"0E9F", X"0AA2", 
		X"FCEC", X"F4DA", X"F105", X"EE6B", X"EC8D", X"EB3C", 
		X"EA75", X"EA27", X"EA51", X"EAF3", X"EC1B", X"EDC9", 
		X"F032", X"F381", X"F8F7", X"08CF", X"0D6C", X"106C", 
		X"1290", X"1413", X"150F", X"158E", X"1596", X"1526", 
		X"143D", X"12CA", X"10C1", X"0DEF", X"09A8", X"FAD2", 
		X"F453", X"F0D8", X"EE69", X"ECA5", X"EB7A", X"EACC", 
		X"EA9B", X"EAE1", X"EBA5", X"ECE7", X"EEC9", X"F158", 
		X"F506", X"FD5D", X"0A60", X"0E3F", X"10E2", X"12C4", 
		X"1412", X"14DA", X"152A", X"1502", X"1462", X"1340", 
		X"1195", X"0F40", X"0BE5", X"0635", X"F708", X"F2B0", 
		X"EFD8", X"EDC9", X"EC61", X"EB7C", X"EB18", X"EB2B", 
		X"EBBA", X"ECC4", X"EE64", X"F0A1", X"F3C9", X"F930", 
		X"0856", X"0CE1", X"0FCD", X"11DE", X"1351", X"143B", 
		X"14A9", X"14A0", X"141F", X"131E", X"1198", X"0F6F", 
		X"0C59", X"0774", X"F83C", X"F383", X"F08A", X"EE68", 
		X"ECF4", X"EC07", X"EB94", X"EB9D", X"EC22", X"ED22", 
		X"EEAA", X"F0E7", X"F3FF", X"F94E", X"0831", X"0CA7", 
		X"0F84", X"1189", X"12EF", X"13D0", X"1434", X"1420", 
		X"1394", X"128B", X"10F3", X"0EB7", X"0B8A", X"05FF", 
		X"F76E", X"F327", X"F06C", X"EE7E", X"ED25", X"EC58", 
		X"EC06", X"EC2D", X"ECCD", X"EDF5", X"EFA5", X"F205", 
		X"F596", X"FCD8", X"09B3", X"0D68", X"0FE8", X"11AD", 
		X"12DC", X"138A", X"13BF", X"137C", X"12BE", X"1180", 
		X"0FAE", X"0D14", X"093D", X"FBB7", X"F550", X"F207", 
		X"EFBB", X"EE28", X"ED21", X"EC97", X"EC89", X"ECF6", 
		X"EDDD", X"EF4A", X"F167", X"F456", X"F91B", X"07B3", 
		X"0C12", X"0ED6", X"10C8", X"121C", X"12EB", X"133F", 
		X"131C", X"127F", X"1165", X"0FBD", X"0D5B", X"09E9", 
		X"017A", X"F650", X"F2D3", X"F06E", X"EECA", X"EDB6", 
		X"ED1F", X"ED04", X"ED63", X"EE3C", X"EF99", X"F1A2", 
		X"F478", X"F90A", X"075B", X"0BB7", X"0E75", X"105D", 
		X"11A9", X"1272", X"12C0", X"1297", X"11F5", X"10D5", 
		X"0F20", X"0CB8", X"0927", X"FC81", X"F5FF", X"F2C6", 
		X"F08B", X"EF07", X"EE0E", X"ED91", X"ED8E", X"EE06", 
		X"EEF8", X"F072", X"F2A2", X"F5BA", X"FB6B", X"0888", 
		X"0C39", X"0EA7", X"1059", X"1177", X"1216", X"123C", 
		X"11ED", X"1123", X"0FD7", X"0DF3", X"0B34", X"06D5", 
		X"F92E", X"F4C8", X"F21E", X"F03D", X"EF01", X"EE47", 
		X"EE05", X"EE3C", X"EEE9", X"F020", X"F1E3", X"F467", 
		X"F873", X"05CE", X"0A93", X"0D5F", X"0F4B", X"109C", 
		X"1165", X"11B6", X"1191", X"10F6", X"0FDE", X"0E32", 
		X"0BD3", X"082B", X"FB6E", X"F60F", X"F317", X"F11B", 
		X"EFC1", X"EEE9", X"EE91", X"EEAD", X"EF43", X"F053", 
		X"F1F0", X"F454", X"F7DF", X"045E", X"09C4", X"0CAB", 
		X"0EA6", X"0FFE", X"10D1", X"112B", X"1110", X"1080", 
		X"0F72", X"0DDA", X"0B8F", X"0807", X"FBB2", X"F650", 
		X"F378", X"F189", X"F035", X"EF6B", X"EF1A", X"EF3F", 
		X"EFD8", X"F0ED", X"F29D", X"F4FE", X"F8AE", X"0583", 
		X"0A07", X"0CAC", X"0E7A", X"0FAF", X"1064", X"10A2", 
		X"106D", X"0FC2", X"0E9A", X"0CE2", X"0A5B", X"0651", 
		X"F9B2", X"F5A3", X"F332", X"F187", X"F068", X"EFCE", 
		X"EFA9", X"EFF8", X"F0BB", X"F209", X"F3E9", X"F6A5", 
		X"FBDF", X"07AD", X"0AFC", X"0D25", X"0E9C", X"0F8B", 
		X"1001", X"1004", X"0F96", X"0EAF", X"0D45", X"0B37", 
		X"0816", X"FD5F", X"F74B", X"F479", X"F296", X"F14B", 
		X"F089", X"F03C", X"F062", X"F0FA", X"F20B", X"F3B5", 
		X"F613", X"F9E4", X"061C", X"09E4", X"0C36", X"0DCA", 
		X"0ED0", X"0F5D", X"0F77", X"0F22", X"0E5A", X"0D0F", 
		X"0B2D", X"0865", X"024D", X"F824", X"F52B", X"F340", 
		X"F1F6", X"F129", X"F0D6", X"F0F2", X"F182", X"F286", 
		X"F413", X"F668", X"FA18", X"05BC", X"0978", X"0BBB", 
		X"0D42", X"0E40", X"0EC5", X"0EDB", X"0E82", X"0DB8", 
		X"0C72", X"0A8B", X"07B8", X"FE62", X"F809", X"F55B", 
		X"F395", X"F261", X"F1B1", X"F171", X"F1A0", X"F23D", 
		X"F350", X"F4FB", X"F761", X"FB94", X"06AB", X"09BE", 
		X"0BB4", X"0D07", X"0DD8", X"0E37", X"0E2A", X"0DB1", 
		X"0CC3", X"0B57", X"0941", X"05E1", X"FAEB", X"F73E", 
		X"F508", X"F394", X"F2A6", X"F22A", X"F21D", X"F27A", 
		X"F34B", X"F494", X"F677", X"F978", X"03D0", X"0810", 
		X"0A5F", X"0BE9", X"0CE8", X"0D74", X"0D94", X"0D4C", 
		X"0C96", X"0B6C", X"09B2", X"070E", X"FE36", X"F8AD", 
		X"F631", X"F496", X"F38A", X"F2EF", X"F2C3", X"F2FE", 
		X"F3A6", X"F4BF", X"F661", X"F8EA", X"FEF1", X"06F6", 
		X"096E", X"0B0A", X"0C18", X"0CB3", X"0CE4", X"0CB1", 
		X"0C14", X"0B0A", X"0979", X"071A", X"0227", X"F96A", 
		X"F6E8", X"F550", X"F445", X"F3A9", X"F379", X"F3AC", 
		X"F449", X"F552", X"F6DE", X"F946", X"FEFF", X"069B", 
		X"08F1", X"0A75", X"0B72", X"0BFF", X"0C29", X"0BF0", 
		X"0B54", X"0A49", X"08BD", X"0666", X"FE64", X"F969", 
		X"F737", X"F5C3", X"F4D9", X"F45A", X"F43D", X"F480", 
		X"F526", X"F63F", X"F7DA", X"FA52", X"0341", X"06DF", 
		X"08D2", X"0A1A", X"0AE8", X"0B50", X"0B59", X"0B05", 
		X"0A50", X"092C", X"077D", X"04CF", X"FBE5", X"F8F0", 
		X"F735", X"F60E", X"F55E", X"F510", X"F51E", X"F587", 
		X"F650", X"F792", X"F967", X"FC9F", X"04FD", X"075B", 
		X"08D5", X"09CA", X"0A58", X"0A89", X"0A62", X"09E1", 
		X"0900", X"07AE", X"05A7", X"0000", X"FA65", X"F86E", 
		X"F732", X"F669", X"F5FF", X"F5EF", X"F634", X"F6D6", 
		X"F7D6", X"F952", X"FBC8", X"03A5", X"0643", X"07C8", 
		X"08C5", X"095B", X"099A", X"0986", X"0920", X"0863", 
		X"073D", X"058A", X"0250", X"FB43", X"F95B", X"F828", 
		X"F763", X"F6FC", X"F6E6", X"F721", X"F7AB", X"F88D", 
		X"F9E9", X"FC02", X"030F", X"0588", X"06EE", X"07D3", 
		X"085B", X"0893", X"087E", X"081F", X"0770", X"0666", 
		X"04D8", X"01AD", X"FBB0", X"FA0C", X"F901", X"F85F", 
		X"F80D", X"F804", X"F843", X"F8C9", X"F99E", X"FAE5", 
		X"FCEE", X"0324", X"050C", X"062B", X"06DF", X"0744", 
		X"0762", X"073F", X"06D9", X"062D", X"052D", X"03AA", 
		X"FE54", X"FBE4", X"FAB0", X"F9ED", X"F97D", X"F951", 
		X"F962", X"F9B0", X"FA3B", X"FB13", X"FC4C", X"FEB8", 
		X"034A", X"0483", X"0542", X"05B3", X"05E5", X"05DF", 
		X"05A4", X"0533", X"0487", X"038F", X"01EB", X"FD8C", 
		X"FC56", X"FBA0", X"FB38", X"FB09", X"FB0C", X"FB3D", 
		X"FB9A", X"FC27", X"FCF4", X"FE29", X"01C0", X"02D0", 
		X"0362", X"03B1", X"03CF", X"03C4", X"0395", X"0344", 
		X"02D2", X"023B", X"016B", X"FF05", X"FE4E", X"FE07", 
		X"FDF7", X"FE13", X"FE55", X"FEBE", X"FF74" );
				
end package sounds;